`ifndef APB_PKT__SV
`define APB_PKT__SV

package apb_pkg;
    import uvm_pkg::*;
    `include "apb_trans.sv"
    `include "apb_sequence.sv"
    `include "apb_sequencer.sv"
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_agent.sv"
    `include "apb_scoreboard.sv"
    `include "apb_coverage.sv"
    `include "apb_env.sv"
endpackage

`endif