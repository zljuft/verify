`ifndef MACROS__VH
`define MACROS__VH

`define AWIDTH 32
`define DWIDTH 32

`endif